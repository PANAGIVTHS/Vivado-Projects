
module FourDigitLEDdriver(reset, clk, appended_byte, append_sig, error, an3, an2, an1, an0, a, b, c, d, e, f, g, dp);
    input clk, reset;
    output an3, an2, an1, an0;
    output wire a, b, c, d, e, f, g, dp;
    wire [3:0] counter;
    wire button_debounced, an3, an2, an1, an0, feedback;
    wire button_ON, enabled, reset_debounced, locked;
    wire [3:0] char;
    input append_sig;
    input error;
    input [7:0] appended_byte;
    
    assign dp = !error;
    
    MMCME2_BASE #(
        .CLKFBOUT_MULT_F(6.0),       // Multiply value for all CLKOUT (2.000-64.000).
        .CLKIN1_PERIOD(10.0),        // Input clock period for 100 MHz clock.
        .CLKOUT0_DIVIDE_F(120.0),    // Divide value for CLKOUT0 to achieve 5 MHz.
        .DIVCLK_DIVIDE(1)            // Divide the input clock by 1.
    )
    MMCME2_BASE_inst (
        .CLKOUT0(new_clk),           // Output: New clock generated by MMCM
        .CLKFBOUT(feedback),         // Output: Feedback clock
        .CLKIN1(clk),                // Input: 100 MHz input clock
        .CLKFBIN(feedback),          // Input: Feedback clock
        .LOCKED(locked)              // Output: Lock signal, high when clock is stable no need to check for this (not that important) + no time
    );

    // if other clock slower then hold to step 
    ConstCounter ConstCounter_inst (.clk(new_clk), .reset(reset), .counter(counter));
    CharacterDecoder CharacterDecoder_inst (.clk(clk), .appended_byte(appended_byte), .append_sig(append_sig), .counter(counter), .char(char), .reset(reset));
    AnodeDecoder AnodeDecoder_inst (.counter(counter), .an0(an0), .an1(an1), .an2(an2), .an3(an3));
    LEDdecoder LEDdecoder_inst (.char(char), .LED({a, b, c, d, e, f, g}));
endmodule
