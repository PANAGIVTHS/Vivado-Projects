
module FRAME7 (
    input clk,
    input reset,
    input read_enable,
    input [1:0] write_enable,
    input reg_enable,
    input [13:0] address,
    output pixel_val
);
   wire [15:0] doa_data;
   wire [15:0] dob_data;      // Unused output for port B
   wire [1:0] dipa_unused;    // Unused parity input for port A
   wire [1:0] dipb_unused;    // Unused parity input for port B
   wire [1:0] dopa_unused;    // Unused parity output for port A
   wire [1:0] dopb_unused;    // Unused parity output for port B

   // RAMB18E1: 18K-bit Configurable Synchronous Block RAM
   //           Artix-7
   // Xilinx HDL Language Template, version 2020.2.
   
   assign dipa_unused = 2'h00;
   assign dipb_unused = 2'h00;
   assign dopa_unused = 2'h00;
   assign dopb_unused = 2'h00;

   RAMB18E1 #(
      .RDADDR_COLLISION_HWCONFIG("DELAYED_WRITE"),
      .SIM_COLLISION_CHECK("ALL"),
      .DOA_REG(0),
      .DOB_REG(0),
      .INIT_00(256'hFFFFFFFE000000000007FFFFFFFFFFFFFFFFFFFE000000000007FFFFFFFFFFFF),
      .INIT_01(256'hFFFFFFF000000000003FFFFFFFFFFFFFFFFFFFFE000000000007FFFFFFFFFFFF),
      .INIT_02(256'hFFFFFFF000000000003FFFFFFFFFFFFFFFFFFFF000000000003FFFFFFFFFFFFF),
      .INIT_03(256'hFFFFFFC00000000000FFFFFFFFFFFFFFFFFFFFC00000000000FFFFFFFFFFFFFF),
      .INIT_04(256'hFFFFFFC00000000000FFFFFFFFFFFFFFFFFFFFC00000000000FFFFFFFFFFFFFF),
      .INIT_05(256'hFFFFFFC00000000000FFFFFFFFFFFFFFFFFFFFC00000000000FFFFFFFFFFFFFF),
      .INIT_06(256'hFFFFFE0000000000003FFFFFFFFFFFFFFFFFFE0000000000003FFFFFFFFFFFFF),
      .INIT_07(256'hFFFFFE0000000000003FFFFFFFFFFFFFFFFFFE0000000000003FFFFFFFFFFFFF),
      .INIT_08(256'hFFFFFE0000000000003FFFFFFFFFFFFFFFFFFE0000000000003FFFFFFFFFFFFF),
      .INIT_09(256'hFFFFF000000000000007FFFFFFFFFFFFFFFFF000000000000007FFFFFFFFFFFF),
      .INIT_0A(256'hFFFFF000000000000007FFFFFFFFFFFFFFFFF000000000000007FFFFFFFFFFFF),
      .INIT_0B(256'hFFFFF000000000000007FFFFFFFFFFFFFFFFF000000000000007FFFFFFFFFFFF),
      .INIT_0C(256'hFFFFF000000000000007FFFFFFFFFFFFFFFFF000000000000007FFFFFFFFFFFF),
      .INIT_0D(256'hFFFFF000000000000007FFFFFFFFFFFFFFFFF000000000000007FFFFFFFFFFFF),
      .INIT_0E(256'hFFFFF000000000000007FFFFFFFFFFFFFFFFF000000000000007FFFFFFFFFFFF),
      .INIT_0F(256'hFFFFC000000000000007FFFFFFFFFFFFFFFFC000000000000007FFFFFFFFFFFF),
      .INIT_10(256'hFFFFC000000000000007FFFFFFFFFFFFFFFFC000000000000007FFFFFFFFFFFF),
      .INIT_11(256'hFFFFC000000000000007FFFFFFFFFFFFFFFFC000000000000007FFFFFFFFFFFF),
      .INIT_12(256'hFFFFC000000000000007FFFFFFFFFFFFFFFFC000000000000007FFFFFFFFFFFF),
      .INIT_13(256'hFFFFC00000000000003FFFFFFFFFFFFFFFFFC000000000000007FFFFFFFFFFFF),
      .INIT_14(256'hFFFFC00000000000003FFFFFFFFFFFFFFFFFC00000000000003FFFFFFFFFFFFF),
      .INIT_15(256'hFFFE000000000001FFFFFFFFFFFFFFFFFFFE000000000001FFFFFFFFFFFFFFFF),
      .INIT_16(256'hFFFE000000000001FFFFFFFFFFFFFFFFFFFE000000000001FFFFFFFFFFFFFFFF),
      .INIT_17(256'hFFFE000000000001FFFFFFFFFFFFFFFFFFFE000000000001FFFFFFFFFFFFFFFF),
      .INIT_18(256'hFFFFC00000000001FFFFFFFFFFFFFFFFFFFFC00000000001FFFFFFFFFFFFFFFF),
      .INIT_19(256'hFFFFC00000000001FFFFFFFFFFFFFFFFFFFFC00000000001FFFFFFFFFFFFFFFF),
      .INIT_1A(256'hFFFFC00000000001FFFFFFFFFFFFFFFFFFFFC00000000001FFFFFFFFFFFFFFFF),
      .INIT_1B(256'hFFFFC00000000007FFFFFFFFFFFFFFFFFFFFC00000000007FFFFFFFFFFFFFFFF),
      .INIT_1C(256'hFFFFC00000000007FFFFFFFFFFFFFFFFFFFFC00000000007FFFFFFFFFFFFFFFF),
      .INIT_1D(256'hFFFFC00000000007FFFFFFFFFFFFFFFFFFFFC00000000007FFFFFFFFFFFFFFFF),
      .INIT_1E(256'hFFFE0E000001C007FFFFFFFFFFFFFFFFFFFE0E000001C007FFFFFFFFFFFFFFFF),
      .INIT_1F(256'hFFFFFE0000000007FFFFFFFFFFFFFFFFFFFE0E000001C007FFFFFFFFFFFFFFFF),
      .INIT_20(256'hFFFFFE0000000007FFFFFFFFFFFFFFFFFFFFFE0000000007FFFFFFFFFFFFFFFF),
      .INIT_21(256'hFFFFFE0000000607FFFFFFFFFFFFFFFFFFFFFE0000000007FFFFFFFFFFFFFFFF),
      .INIT_22(256'hFFFFFE0000000607FFFFFFFFFFFFFFFFFFFFFE0000000607FFFFFFFFFFFFFFFF),
      .INIT_23(256'hFFFFFE0000000007FFFFFFFFFFFFFFFFFFFFFE0000000007FFFFFFFFFFFFFFFF),
      .INIT_24(256'hFFFFF0000000003FFFFFFFFFFFFFFFFFFFFFFE0000000007FFFFFFFFFFFFFFFF),
      .INIT_25(256'hFFFFF0000000003FFFFFFFFFFFFFFFFFFFFFF0000000003FFFFFFFFFFFFFFFFF),
      .INIT_26(256'hFFFFF0000000003FFFFFFFFFFFFFFFFFFFFFF0000000003FFFFFFFFFFFFFFFFF),
      .INIT_27(256'hFFFFC0000000003FFFFFC0003FFFFFFFFFFFF0000000003FFFFFFFFFFFFFFFFF),
      .INIT_28(256'hFFFFC0000000003FFFFFC0003FFFFFFFFFFFC0000000003FFFFFC0003FFFFFFF),
      .INIT_29(256'hFFFFC0000000003FFFFFC0003FFFFFFFFFFFC0000000003FFFFFC0003FFFFFFF),
      .INIT_2A(256'hFFFFF0000000003FFFFF000007FFFFFFFFFFC0000000003FFFFFC0003FFFFFFF),
      .INIT_2B(256'hFFFFF0000000003FFFFF000007FFFFFFFFFFF0000000003FFFFF000007FFFFFF),
      .INIT_2C(256'hFFFFF0000000003FFFF8000007FFFFFFFFFFF0000000003FFFF8000007FFFFFF),
      .INIT_2D(256'hFFFFC0000000003FFF00000007FFFFFFFFFFF0000000003FFFF8000007FFFFFF),
      .INIT_2E(256'hFFFFC0000000003FFF00000007FFFFFFFFFFC0000000003FFF00000007FFFFFF),
      .INIT_2F(256'hFFFFC0000000003FFF00000007FFFFFFFFFFC0000000003FFF00000007FFFFFF),
      .INIT_A(18'h00000),
      .INIT_B(18'h00000),
      .INIT_FILE("NONE"),
      .RAM_MODE("TDP"),
      .READ_WIDTH_A(1), 
      .READ_WIDTH_B(0), 
      .WRITE_WIDTH_A(0), 
      .WRITE_WIDTH_B(0), 
      .RSTREG_PRIORITY_A("RSTREG"),
      .RSTREG_PRIORITY_B("RSTREG"),
      .SRVAL_A(18'h00000),
      .SRVAL_B(18'h00000),
      .SIM_DEVICE("7SERIES"),
      .WRITE_MODE_A("WRITE_FIRST"),
      .WRITE_MODE_B("WRITE_FIRST")
   )
   RAMB18E1_inst (
      // Port A
      .DOADO(doa_data),                   // 16-bit output: A port data/LSB data
      .DOPADOP(dopa_unused),              // 2-bit output: A port parity data
      .ADDRARDADDR(address),      // 15-bit input: A port address (with MSB padding)
      .CLKARDCLK(clk),                    // 1-bit input: A port clock/Read clock
      .ENARDEN(read_enable),              // 1-bit input: A port enable/Read enable
      .REGCEAREGCE(reg_enable),           // 1-bit input: A port register enable/Register enable
      .RSTRAMARSTRAM(reset),              // 1-bit input: A port set/reset
      .RSTREGARSTREG(reset),              // 1-bit input: A port register set/reset
      .DIADI(16'h0000),                   // 16-bit input: A port data input
      .DIPADIP(dipa_unused),              // 2-bit input: A port parity input
      .WEA(write_enable),                 // 2-bit input: A port write enable

      // Port B (Unused)
      .DOBDO(dob_data),                   // 16-bit output: B port data
      .DOPBDOP(dopb_unused),              // 2-bit output: B port parity data
      .ADDRBWRADDR(14'b0),             // 15-bit input: B port address
      .CLKBWRCLK(1'b0),                   // 1-bit input: B port clock
      .ENBWREN(1'b0),                     // 1-bit input: B port enable
      .REGCEB(1'b0),                      // 1-bit input: B port register enable
      .RSTRAMB(1'b0),                     // 1-bit input: B port set/reset
      .RSTREGB(1'b0),                     // 1-bit input: B port register set/reset
      .DIBDI(16'h0000),                   // 16-bit input: B port data input
      .DIPBDIP(dipb_unused),              // 2-bit input: B port parity input
      .WEBWE(4'b0000)                     // 4-bit input: B port write enable
   );

   assign pixel_val = doa_data[0];

endmodule
