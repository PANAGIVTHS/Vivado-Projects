
module FRAME3 (
    input clk,
    input reset,
    input read_enable,
    input [1:0] write_enable,
    input reg_enable,
    input [13:0] address,
    output pixel_val
);
   wire [15:0] doa_data;
   wire [15:0] dob_data;      // Unused output for port B
   wire [1:0] dipa_unused;    // Unused parity input for port A
   wire [1:0] dipb_unused;    // Unused parity input for port B
   wire [1:0] dopa_unused;    // Unused parity output for port A
   wire [1:0] dopb_unused;    // Unused parity output for port B

   // RAMB18E1: 18K-bit Configurable Synchronous Block RAM
   //           Artix-7
   // Xilinx HDL Language Template, version 2020.2.
   
   assign dipa_unused = 2'h00;
   assign dipb_unused = 2'h00;
   assign dopa_unused = 2'h00;
   assign dopb_unused = 2'h00;

   RAMB18E1 #(
      .RDADDR_COLLISION_HWCONFIG("DELAYED_WRITE"),
      .SIM_COLLISION_CHECK("ALL"),
      .DOA_REG(0),
      .DOB_REG(0),
      .INIT_00(256'hFFFFFFFFFFF800000007FFFFFFFFFFFFFFFFFFFFFFF800000007FFFFFFFFFFFF),
      .INIT_01(256'hFFFFFFFFFFF800000007FFFFFFFFFFFFFFFFFFFFFFF800000007FFFFFFFFFFFF),
      .INIT_02(256'hFFFFFFFFFFF800000007FFFFFFFFFFFFFFFFFFFFFFF800000007FFFFFFFFFFFF),
      .INIT_03(256'hFFFFFFFFFFF800000007FFFFFFFFFFFFFFFFFFFFFFF800000007FFFFFFFFFFFF),
      .INIT_04(256'hFFFFFFFFFFF800000007FFFFFFFFFFFFFFFFFFFFFFF800000007FFFFFFFFFFFF),
      .INIT_05(256'hFFFFFFFFFFFF0000001FFFFFFFFFFFFFFFFFFFFFFFF800000007FFFFFFFFFFFF),
      .INIT_06(256'hFFFFFFFFFFFF0000001FFFFFFFFFFFFFFFFFFFFFFFFF0000001FFFFFFFFFFFFF),
      .INIT_07(256'hFFFFFFFFFFFF0000001FFFFFFFFFFFFFFFFFFFFFFFFF0000001FFFFFFFFFFFFF),
      .INIT_08(256'hFFFFFFFFFFFF0000001FFFFFFFFFFFFFFFFFFFFFFFFF0000001FFFFFFFFFFFFF),
      .INIT_09(256'hFFFFFFFFFFFF0000001FFFFFFFFFFFFFFFFFFFFFFFFF0000001FFFFFFFFFFFFF),
      .INIT_0A(256'hFFFFFFFFFFFF000000FFFFFFFFFFFFFFFFFFFFFFFFFF000000FFFFFFFFFFFFFF),
      .INIT_0B(256'hFFFFFFFFFFFF000007FFFFFFFFFFFFFFFFFFFFFFFFFF000000FFFFFFFFFFFFFF),
      .INIT_0C(256'hFFFFFFFFFFFF000007FFFFFFFFFFFFFFFFFFFFFFFFFF000007FFFFFFFFFFFFFF),
      .INIT_0D(256'hFFFFFFFFFFFF000007FFFFFFFFFFFFFFFFFFFFFFFFFF000007FFFFFFFFFFFFFF),
      .INIT_0E(256'hFFFFFFFFFFFF000007FFFFFFFFFFFFFFFFFFFFFFFFFF000007FFFFFFFFFFFFFF),
      .INIT_0F(256'hFFFFFFFFFFFF000007FFFFFFFFFFFFFFFFFFFFFFFFFF000007FFFFFFFFFFFFFF),
      .INIT_10(256'hFFFFFFFFFFFF000000FFFFFFFFFFFFFFFFFFFFFFFFFF000007FFFFFFFFFFFFFF),
      .INIT_11(256'hFFFFFFFFFFFF000000FFFFFFFFFFFFFFFFFFFFFFFFFF000000FFFFFFFFFFFFFF),
      .INIT_12(256'hFFFFFFFFFFFF0000001FFFFFFFFFFFFFFFFFFFFFFFFF0000001FFFFFFFFFFFFF),
      .INIT_13(256'hFFFFFFFFFFFF0000001FFFFFFFFFFFFFFFFFFFFFFFFF0000001FFFFFFFFFFFFF),
      .INIT_14(256'hFFFFFFFFFFFF0000001FFFFFFFFFFFFFFFFFFFFFFFFF0000001FFFFFFFFFFFFF),
      .INIT_15(256'hFFFFFFFFFFFF0000001FFFFFFFFFFFFFFFFFFFFFFFFF0000001FFFFFFFFFFFFF),
      .INIT_16(256'hFFFFFFFFFFFF0000001FFFFFFFFFFFFFFFFFFFFFFFFF0000001FFFFFFFFFFFFF),
      .INIT_17(256'hFFFFFFFFFFFF0000001FFFFFFFFFFFFFFFFFFFFFFFFF0000001FFFFFFFFFFFFF),
      .INIT_18(256'hFFFFFFFFFFF800000007FFFFFFFFFFFFFFFFFFFFFFF800000007FFFFFFFFFFFF),
      .INIT_19(256'hFFFFFFFFFFF800000007FFFFFFFFFFFFFFFFFFFFFFF800000007FFFFFFFFFFFF),
      .INIT_1A(256'hFFFFFFFFFFF800000007FFFFFFFFFFFFFFFFFFFFFFF800000007FFFFFFFFFFFF),
      .INIT_1B(256'hFFFFFFFFFFF800000000FFFFFFFFFFFFFFFFFFFFFFF800000000FFFFFFFFFFFF),
      .INIT_1C(256'hFFFFFFFFFFF800000000FFFFFFFFFFFFFFFFFFFFFFF800000000FFFFFFFFFFFF),
      .INIT_1D(256'hFFFFFFFFFFF800000000FFFFFFFFFFFFFFFFFFFFFFF800000000FFFFFFFFFFFF),
      .INIT_1E(256'hFFFFFFFFFFC03F0000001FFFFFFFFFFFFFFFFFFFFFC03F0000001FFFFFFFFFFF),
      .INIT_1F(256'hFFFFFFFFFFC03F0000001FFFFFFFFFFFFFFFFFFFFFC03F0000001FFFFFFFFFFF),
      .INIT_20(256'hFFFFFFFFFFC03F0000001FFFFFFFFFFFFFFFFFFFFFC03F0000001FFFFFFFFFFF),
      .INIT_21(256'hFFFFFFFFFF003F00000007FFFFFFFFFFFFFFFFFFFF003F00000007FFFFFFFFFF),
      .INIT_22(256'hFFFFFFFFFF003F00000007FFFFFFFFFFFFFFFFFFFF003F00000007FFFFFFFFFF),
      .INIT_23(256'hFFFFFFFFFF003F00000007FFFFFFFFFFFFFFFFFFFF003F00000007FFFFFFFFFF),
      .INIT_24(256'hFFFFFFFFF8003800000007FFFFFFFFFFFFFFFFFFFF003F00000007FFFFFFFFFF),
      .INIT_25(256'hFFFFFFFFF8003800000007FFFFFFFFFFFFFFFFFFF8003800000007FFFFFFFFFF),
      .INIT_26(256'hFFFFFFFFF8000000000007FFFFFFFFFFFFFFFFFFF8000000000007FFFFFFFFFF),
      .INIT_27(256'hFFFFFFFFF8000000000007FFFFFFFFFFFFFFFFFFF8000000000007FFFFFFFFFF),
      .INIT_28(256'hFFFFFFFFF8000000000007FFFFFFFFFFFFFFFFFFF8000000000007FFFFFFFFFF),
      .INIT_29(256'hFFFFFFFFF8000000000007FFFFFFFFFFFFFFFFFFF8000000000007FFFFFFFFFF),
      .INIT_2A(256'hFFFFFFFFF800000000001FFFFFFFFFFFFFFFFFFFF8000000000007FFFFFFFFFF),
      .INIT_2B(256'hFFFFFFFFF800000000001FFFFFFFFFFFFFFFFFFFF800000000001FFFFFFFFFFF),
      .INIT_2C(256'hFFFFFFFFF800000000001FFFFFFFFFFFFFFFFFFFF800000000001FFFFFFFFFFF),
      .INIT_2D(256'hFFFFFFFFF83F00000000FFFFFFFFFFFFFFFFFFFFF800000000001FFFFFFFFFFF),
      .INIT_2E(256'hFFFFFFFFF83F00000000FFFFFFFFFFFFFFFFFFFFF83F00000000FFFFFFFFFFFF),
      .INIT_2F(256'hFFFFFFFFF83F00000000FFFFFFFFFFFFFFFFFFFFF83F00000000FFFFFFFFFFFF),
      .INIT_A(18'h00000),
      .INIT_B(18'h00000),
      .INIT_FILE("NONE"),
      .RAM_MODE("TDP"),
      .READ_WIDTH_A(1), 
      .READ_WIDTH_B(0), 
      .WRITE_WIDTH_A(0), 
      .WRITE_WIDTH_B(0), 
      .RSTREG_PRIORITY_A("RSTREG"),
      .RSTREG_PRIORITY_B("RSTREG"),
      .SRVAL_A(18'h00000),
      .SRVAL_B(18'h00000),
      .SIM_DEVICE("7SERIES"),
      .WRITE_MODE_A("WRITE_FIRST"),
      .WRITE_MODE_B("WRITE_FIRST")
   )
   RAMB18E1_inst (
      // Port A
      .DOADO(doa_data),                   // 16-bit output: A port data/LSB data
      .DOPADOP(dopa_unused),              // 2-bit output: A port parity data
      .ADDRARDADDR(address),      // 15-bit input: A port address (with MSB padding)
      .CLKARDCLK(clk),                    // 1-bit input: A port clock/Read clock
      .ENARDEN(read_enable),              // 1-bit input: A port enable/Read enable
      .REGCEAREGCE(reg_enable),           // 1-bit input: A port register enable/Register enable
      .RSTRAMARSTRAM(reset),              // 1-bit input: A port set/reset
      .RSTREGARSTREG(reset),              // 1-bit input: A port register set/reset
      .DIADI(16'h0000),                   // 16-bit input: A port data input
      .DIPADIP(dipa_unused),              // 2-bit input: A port parity input
      .WEA(write_enable),                 // 2-bit input: A port write enable

      // Port B (Unused)
      .DOBDO(dob_data),                   // 16-bit output: B port data
      .DOPBDOP(dopb_unused),              // 2-bit output: B port parity data
      .ADDRBWRADDR(14'h0000),             // 15-bit input: B port address
      .CLKBWRCLK(1'b0),                   // 1-bit input: B port clock
      .ENBWREN(1'b0),                     // 1-bit input: B port enable
      .REGCEB(1'b0),                      // 1-bit input: B port register enable
      .RSTRAMB(1'b0),                     // 1-bit input: B port set/reset
      .RSTREGB(1'b0),                     // 1-bit input: B port register set/reset
      .DIBDI(16'h0000),                   // 16-bit input: B port data input
      .DIPBDIP(dipb_unused),              // 2-bit input: B port parity input
      .WEBWE(4'b0000)                     // 4-bit input: B port write enable
   );

   assign pixel_val = doa_data[0];

endmodule
