
module FRAME1 (
    input clk,
    input reset,
    input read_enable,
    input [1:0] write_enable,
    input reg_enable,
    input [13:0] address,
    output pixel_val
);
   wire [15:0] doa_data;
   wire [15:0] dob_data;      // Unused output for port B
   wire [1:0] dipa_unused;    // Unused parity input for port A
   wire [1:0] dipb_unused;    // Unused parity input for port B
   wire [1:0] dopa_unused;    // Unused parity output for port A
   wire [1:0] dopb_unused;    // Unused parity output for port B

   // RAMB18E1: 18K-bit Configurable Synchronous Block RAM
   //           Artix-7
   // Xilinx HDL Language Template, version 2020.2.
   
   assign dipa_unused = 2'h00;
   assign dipb_unused = 2'h00;
   assign dopa_unused = 2'h00;
   assign dopb_unused = 2'h00;

   RAMB18E1 #(
      .RDADDR_COLLISION_HWCONFIG("DELAYED_WRITE"),
      .SIM_COLLISION_CHECK("ALL"),
      .DOA_REG(0),
      .DOB_REG(0),
      .INIT_00(256'hFFFFFFFFFFFF00000000000000000000FFFFFFFFFFFF00000000000000000000),
      .INIT_01(256'hFFFFFFFFFFFF00000000000000000000FFFFFFFFFFFF00000000000000000000),
      .INIT_02(256'hFFFFFFFFFFFF00000000000000000000FFFFFFFFFFFF00000000000000000000),
      .INIT_03(256'hFFFFFFFFFFFFC0000000000000000000FFFFFFFFFFFFC0000000000000000000),
      .INIT_04(256'hFFFFFFFFFFFFF0000000000000000000FFFFFFFFFFFFC0000000000000000000),
      .INIT_05(256'hFFFFFFFFFFFFF0000000000000000000FFFFFFFFFFFFF0000000000000000000),
      .INIT_06(256'hFFFFFFFFFFFFFC000000000000000000FFFFFFFFFFFFFC000000000000000000),
      .INIT_07(256'hFFFFFFFFFFFFFC000000000000000000FFFFFFFFFFFFFC000000000000000000),
      .INIT_08(256'hFFFFFFFFFFFFFC000000000000000000FFFFFFFFFFFFFC000000000000000000),
      .INIT_09(256'hFFFFFFFFFFFFFF000000000000000000FFFFFFFFFFFFFF000000000000000000),
      .INIT_0A(256'hFFFFFFFFFFFFFF000000000000000000FFFFFFFFFFFFFF000000000000000000),
      .INIT_0B(256'hFFFFFFFFFFFFFF000000000000000000FFFFFFFFFFFFFF000000000000000000),
      .INIT_0C(256'hFFFFFFFFFFFFFF000000000000000000FFFFFFFFFFFFFF000000000000000000),
      .INIT_0D(256'hFFFFFFFFFFFFFF000000000000000000FFFFFFFFFFFFFF000000000000000000),
      .INIT_0E(256'hFFFFFFFFFFFFFF000000000000000000FFFFFFFFFFFFFF000000000000000000),
      .INIT_0F(256'hFFFFFFFFFFFFFC000000000000000000FFFFFFFFFFFFFC000000000000000000),
      .INIT_10(256'hFFFFFFFFFFFFF0000000000000000000FFFFFFFFFFFFFC000000000000000000),
      .INIT_11(256'hFFFFFFFFFFFFF0000000000000000000FFFFFFFFFFFFF0000000000000000000),
      .INIT_12(256'hFFFFFFFFFFFF00000000000000000000FFFFFFFFFFFF00000000000000000000),
      .INIT_13(256'hFFFFFFFFFFFF00000000000000000000FFFFFFFFFFFF00000000000000000000),
      .INIT_14(256'hFFFFFFFFFFFF00000000000000000000FFFFFFFFFFFF00000000000000000000),
      .INIT_15(256'hFFFFFFFFFFFFC0000000000000000000FFFFFFFFFFFFC0000000000000000000),
      .INIT_16(256'hFFFFFFFFFFFF00000000000000000000FFFFFFFFFFFFC0000000000000000000),
      .INIT_17(256'hFFFFFFFFFFFF00000000000000000000FFFFFFFFFFFF00000000000000000000),
      .INIT_18(256'hFFFFFFFFFFF000000000000000000000FFFFFFFFFFF000000000000000000000),
      .INIT_19(256'hFFFFFFFFFFC000000000000000000000FFFFFFFFFFF000000000000000000000),
      .INIT_1A(256'hFFFFFFFFFFC000000000000000000000FFFFFFFFFFC000000000000000000000),
      .INIT_1B(256'hFFFFFFFFFC0000000000000000000000FFFFFFFFFC0000000000000000000000),
      .INIT_1C(256'hFFFFFFFFFC0000000000000000000000FFFFFFFFFC0000000000000000000000),
      .INIT_1D(256'hFFFFFFFFFC0000000000000000000000FFFFFFFFFC0000000000000000000000),
      .INIT_1E(256'hFFFFFFFFF00000000000000000000000FFFFFFFFF00000000000000000000000),
      .INIT_1F(256'hFFFFFFFFF00000000000000000000000FFFFFFFFF00000000000000000000000),
      .INIT_20(256'hFFFFFFFFF00000000000000000000000FFFFFFFFF00000000000000000000000),
      .INIT_21(256'hFFFFFFFFC00000000000000000000000FFFFFFFFC00000000000000000000000),
      .INIT_22(256'hFFFFFFFFC00000000000000000000000FFFFFFFFC00000000000000000000000),
      .INIT_23(256'hFFFFFFFFC00000000000000000000000FFFFFFFFC00000000000000000000000),
      .INIT_24(256'hFFFFFFFF000000000000000000000000FFFFFFFF000000000000000000000000),
      .INIT_25(256'hFFFFFFFF000000000000000000000000FFFFFFFF000000000000000000000000),
      .INIT_26(256'hFFFFFFFF000000000000000000000000FFFFFFFF000000000000000000000000),
      .INIT_27(256'hFFFFFFFF000000000000000000000000FFFFFFFF000000000000000000000000),
      .INIT_28(256'hFFFFFFFF000000000000000000000000FFFFFFFF000000000000000000000000),
      .INIT_29(256'hFFFFFFFF000000000000000000000000FFFFFFFF000000000000000000000000),
      .INIT_2A(256'hFFFFFFFF000000000000000000000000FFFFFFFF000000000000000000000000),
      .INIT_2B(256'hFFFFFFFF000000000000000000000000FFFFFFFF000000000000000000000000),
      .INIT_2C(256'hFFFFFFFF000000000000000000000000FFFFFFFF000000000000000000000000),
      .INIT_2D(256'hFFFFFFFC000000000000000000000000FFFFFFFC000000000000000000000000),
      .INIT_2E(256'hFFFFFFFC000000000000000000000000FFFFFFFC000000000000000000000000),
      .INIT_2F(256'hFFFFFFFC000000000000000000000000FFFFFFFC000000000000000000000000),
      .INIT_A(18'h00000),
      .INIT_B(18'h00000),
      .INIT_FILE("NONE"),
      .RAM_MODE("TDP"),
      .READ_WIDTH_A(1), 
      .READ_WIDTH_B(0), 
      .WRITE_WIDTH_A(0), 
      .WRITE_WIDTH_B(0), 
      .RSTREG_PRIORITY_A("RSTREG"),
      .RSTREG_PRIORITY_B("RSTREG"),
      .SRVAL_A(18'h00000),
      .SRVAL_B(18'h00000),
      .SIM_DEVICE("7SERIES"),
      .WRITE_MODE_A("WRITE_FIRST"),
      .WRITE_MODE_B("WRITE_FIRST")
   )
   RAMB18E1_inst (
      // Port A
      .DOADO(doa_data),                   // 16-bit output: A port data/LSB data
      .DOPADOP(dopa_unused),              // 2-bit output: A port parity data
      .ADDRARDADDR(address),      // 15-bit input: A port address (with MSB padding)
      .CLKARDCLK(clk),                    // 1-bit input: A port clock/Read clock
      .ENARDEN(read_enable),              // 1-bit input: A port enable/Read enable
      .REGCEAREGCE(reg_enable),           // 1-bit input: A port register enable/Register enable
      .RSTRAMARSTRAM(reset),              // 1-bit input: A port set/reset
      .RSTREGARSTREG(reset),              // 1-bit input: A port register set/reset
      .DIADI(16'h0000),                   // 16-bit input: A port data input
      .DIPADIP(dipa_unused),              // 2-bit input: A port parity input
      .WEA(write_enable),                 // 2-bit input: A port write enable

      // Port B (Unused)
      .DOBDO(dob_data),                   // 16-bit output: B port data
      .DOPBDOP(dopb_unused),              // 2-bit output: B port parity data
      .ADDRBWRADDR(14'b0),             // 15-bit input: B port address
      .CLKBWRCLK(1'b0),                   // 1-bit input: B port clock
      .ENBWREN(1'b0),                     // 1-bit input: B port enable
      .REGCEB(1'b0),                      // 1-bit input: B port register enable
      .RSTRAMB(1'b0),                     // 1-bit input: B port set/reset
      .RSTREGB(1'b0),                     // 1-bit input: B port register set/reset
      .DIBDI(16'h0000),                   // 16-bit input: B port data input
      .DIPBDIP(dipb_unused),              // 2-bit input: B port parity input
      .WEBWE(4'b0000)                     // 4-bit input: B port write enable
   );

   assign pixel_val = doa_data[0];

endmodule
