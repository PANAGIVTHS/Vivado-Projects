
module FRAME8 (
    input clk,
    input reset,
    input read_enable,
    input [1:0] write_enable,
    input reg_enable,
    input [13:0] address,
    output pixel_val
);
   wire [15:0] doa_data;
   wire [15:0] dob_data;      // Unused output for port B
   wire [1:0] dipa_unused;    // Unused parity input for port A
   wire [1:0] dipb_unused;    // Unused parity input for port B
   wire [1:0] dopa_unused;    // Unused parity output for port A
   wire [1:0] dopb_unused;    // Unused parity output for port B

   // RAMB18E1: 18K-bit Configurable Synchronous Block RAM
   //           Artix-7
   // Xilinx HDL Language Template, version 2020.2.
   
   assign dipa_unused = 2'h00;
   assign dipb_unused = 2'h00;
   assign dopa_unused = 2'h00;
   assign dopb_unused = 2'h00;

   RAMB18E1 #(
      .RDADDR_COLLISION_HWCONFIG("DELAYED_WRITE"),
      .SIM_COLLISION_CHECK("ALL"),
      .DOA_REG(0),
      .DOB_REG(0),
      .INIT_00(256'hFFFFFFFFF8000000000000FFFFFFFFFFFFFFFFFFF8000000000000FFFFFFFFFF),
      .INIT_01(256'hFFFFFFFFF8000000000000FFFFFFFFFFFFFFFFFFF8000000000000FFFFFFFFFF),
      .INIT_02(256'hFFFFFFFFC0000000000000FFFFFFFFFFFFFFFFFFF8000000000000FFFFFFFFFF),
      .INIT_03(256'hFFFFFFFFC0000000000000FFFFFFFFFFFFFFFFFFC0000000000000FFFFFFFFFF),
      .INIT_04(256'hFFFFFFFE00000000000000FFFFFFFFFFFFFFFFFE00000000000000FFFFFFFFFF),
      .INIT_05(256'hFFFFFFF800000000000007FFFFFFFFFFFFFFFFFE00000000000000FFFFFFFFFF),
      .INIT_06(256'hFFFFFFF800000000000007FFFFFFFFFFFFFFFFF800000000000007FFFFFFFFFF),
      .INIT_07(256'hFFFFFFF80000000000001FFFFFFFFFFFFFFFFFF80000000000001FFFFFFFFFFF),
      .INIT_08(256'hFFFFFFC0000000000007FFFFFFFFFFFFFFFFFFF80000000000001FFFFFFFFFFF),
      .INIT_09(256'hFFFFFFC0000000000007FFFFFFFFFFFFFFFFFFC0000000000007FFFFFFFFFFFF),
      .INIT_0A(256'hFFFFFFC0000000000007FFFFFFFFFFFFFFFFFFC0000000000007FFFFFFFFFFFF),
      .INIT_0B(256'hFFFFFE00000000000000FFFFFFFFFFFFFFFFFFC0000000000007FFFFFFFFFFFF),
      .INIT_0C(256'hFFFFFE00000000000000FFFFFFFFFFFFFFFFFE00000000000000FFFFFFFFFFFF),
      .INIT_0D(256'hFFFFFE00000000000000FFFFFFFFFFFFFFFFFE00000000000000FFFFFFFFFFFF),
      .INIT_0E(256'hFFFFFE00000000000000FFFFFFFFFFFFFFFFFE00000000000000FFFFFFFFFFFF),
      .INIT_0F(256'hFFFFFE00000000000000FFFFFFFFFFFFFFFFFE00000000000000FFFFFFFFFFFF),
      .INIT_10(256'hFFFFFE00000000000000FFFFFFFFFFFFFFFFFE00000000000000FFFFFFFFFFFF),
      .INIT_11(256'hFFFFF800000000000000FFFFFFFFFFFFFFFFFE00000000000000FFFFFFFFFFFF),
      .INIT_12(256'hFFFFF800000000000000FFFFFFFFFFFFFFFFF800000000000000FFFFFFFFFFFF),
      .INIT_13(256'hFFFFF800000000000000FFFFFFFFFFFFFFFFF800000000000000FFFFFFFFFFFF),
      .INIT_14(256'hFFFFF800000000000000FFFFFFFFFFFFFFFFF800000000000000FFFFFFFFFFFF),
      .INIT_15(256'hFFFFF800000000000000FFFFFFFFFFFFFFFFF800000000000000FFFFFFFFFFFF),
      .INIT_16(256'hFFFFF800000000000007FFFFFFFFFFFFFFFFF800000000000000FFFFFFFFFFFF),
      .INIT_17(256'hFFFFF800000000000007FFFFFFFFFFFFFFFFF800000000000007FFFFFFFFFFFF),
      .INIT_18(256'hFFFFC0000000000007FFFFFFFFFFFFFFFFFFC0000000000007FFFFFFFFFFFFFF),
      .INIT_19(256'hFFFFC0000000000007FFFFFFFFFFFFFFFFFFC0000000000007FFFFFFFFFFFFFF),
      .INIT_1A(256'hFFFFC0000000000007FFFFFFFFFFFFFFFFFFC0000000000007FFFFFFFFFFFFFF),
      .INIT_1B(256'hFFFFC000000000001FFFFFFFFFFFFFFFFFFFC000000000001FFFFFFFFFFFFFFF),
      .INIT_1C(256'hFFFFC000000000001FFFFFFFFFFFFFFFFFFFC000000000001FFFFFFFFFFFFFFF),
      .INIT_1D(256'hFFFFC000000000001FFFFFFFFFFFFFFFFFFFC000000000001FFFFFFFFFFFFFFF),
      .INIT_1E(256'hFFFFC0000007C0F81FFFFFFFFFFFFFFFFFFFC0000007C0F81FFFFFFFFFFFFFFF),
      .INIT_1F(256'hFFFFC0000007C0F81FFFFFFFFFFFFFFFFFFFC0000007C0F81FFFFFFFFFFFFFFF),
      .INIT_20(256'hFFFFC0000007C0F81FFFFFFFFFFFFFFFFFFFC0000007C0F81FFFFFFFFFFFFFFF),
      .INIT_21(256'hFFFFF8000000C0F81FFFFFFFFFFFFFFFFFFFF8000000C0F81FFFFFFFFFFFFFFF),
      .INIT_22(256'hFFFFF800000000F81FFFFFFFFFFFFFFFFFFFF8000000C0F81FFFFFFFFFFFFFFF),
      .INIT_23(256'hFFFFF800000000F81FFFFFFFFFFFFFFFFFFFF800000000F81FFFFFFFFFFFFFFF),
      .INIT_24(256'hFFFFC000000007F81FFFFFFFFFFFFFFFFFFFC000000007F81FFFFFFFFFFFFFFF),
      .INIT_25(256'hFFFE0000000007F81FFFFFFFFFFFFFFFFFFFC000000007F81FFFFFFFFFFFFFFF),
      .INIT_26(256'hFFFE0000000007F81FFFFFFFFFFFFFFFFFFE0000000007F81FFFFFFFFFFFFFFF),
      .INIT_27(256'hFFF80000000007F8FFFFFFFFFFFFFFFFFFF80000000007F8FFFFFFFFFFFFFFFF),
      .INIT_28(256'hFFF80000000007FFFFFFFFFFFFFFFFFFFFF80000000007F8FFFFFFFFFFFFFFFF),
      .INIT_29(256'hFFF80000000007FFFFFFFFFFFFFFFFFFFFF80000000007FFFFFFFFFFFFFFFFFF),
      .INIT_2A(256'hFFC00000000000FFFFFFFFFFFFFFFFFFFFC00000000000FFFFFFFFFFFFFFFFFF),
      .INIT_2B(256'hFFC00000000000FFFFFFFFFFFFFFFFFFFFC00000000000FFFFFFFFFFFFFFFFFF),
      .INIT_2C(256'hFFC00000000000FFFFFFFFFFFFFFFFFFFFC00000000000FFFFFFFFFFFFFFFFFF),
      .INIT_2D(256'hFE000000000007FFFFFFFFFFFFFFFFFFFE000000000007FFFFFFFFFFFFFFFFFF),
      .INIT_2E(256'hFE000000000007FFFFFFFFFFFFFFFFFFFE000000000007FFFFFFFFFFFFFFFFFF),
      .INIT_2F(256'hFE000000000007FFFFFFFFFFFFFFFFFFFE000000000007FFFFFFFFFFFFFFFFFF),
      .INIT_A(18'h00000),
      .INIT_B(18'h00000),
      .INIT_FILE("NONE"),
      .RAM_MODE("TDP"),
      .READ_WIDTH_A(1), 
      .READ_WIDTH_B(0), 
      .WRITE_WIDTH_A(0), 
      .WRITE_WIDTH_B(0), 
      .RSTREG_PRIORITY_A("RSTREG"),
      .RSTREG_PRIORITY_B("RSTREG"),
      .SRVAL_A(18'h00000),
      .SRVAL_B(18'h00000),
      .SIM_DEVICE("7SERIES"),
      .WRITE_MODE_A("WRITE_FIRST"),
      .WRITE_MODE_B("WRITE_FIRST")
   )
   RAMB18E1_inst (
      // Port A
      .DOADO(doa_data),                   // 16-bit output: A port data/LSB data
      .DOPADOP(dopa_unused),              // 2-bit output: A port parity data
      .ADDRARDADDR(address),      // 15-bit input: A port address (with MSB padding)
      .CLKARDCLK(clk),                    // 1-bit input: A port clock/Read clock
      .ENARDEN(read_enable),              // 1-bit input: A port enable/Read enable
      .REGCEAREGCE(reg_enable),           // 1-bit input: A port register enable/Register enable
      .RSTRAMARSTRAM(reset),              // 1-bit input: A port set/reset
      .RSTREGARSTREG(reset),              // 1-bit input: A port register set/reset
      .DIADI(16'h0000),                   // 16-bit input: A port data input
      .DIPADIP(dipa_unused),              // 2-bit input: A port parity input
      .WEA(write_enable),                 // 2-bit input: A port write enable

      // Port B (Unused)
      .DOBDO(dob_data),                   // 16-bit output: B port data
      .DOPBDOP(dopb_unused),              // 2-bit output: B port parity data
      .ADDRBWRADDR(14'b0),             // 15-bit input: B port address
      .CLKBWRCLK(1'b0),                   // 1-bit input: B port clock
      .ENBWREN(1'b0),                     // 1-bit input: B port enable
      .REGCEB(1'b0),                      // 1-bit input: B port register enable
      .RSTRAMB(1'b0),                     // 1-bit input: B port set/reset
      .RSTREGB(1'b0),                     // 1-bit input: B port register set/reset
      .DIBDI(16'h0000),                   // 16-bit input: B port data input
      .DIPBDIP(dipb_unused),              // 2-bit input: B port parity input
      .WEBWE(4'b0000)                     // 4-bit input: B port write enable
   );

   assign pixel_val = doa_data[0];

endmodule
